----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:49:06 02/13/2026 
-- Design Name: 
-- Module Name:    LAB_1A - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LAB_1A is
    Port ( color_in : in  STD_LOGIC_VECTOR (11 downto 0);
           color_out : out  STD_LOGIC_VECTOR (11 downto 0));
end LAB_1A;

architecture Behavioral of LAB_1A is

begin


end Behavioral;

